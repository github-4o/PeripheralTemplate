library ieee;
use ieee.std_logic_1164.all;


package platform is

    constant cAsync_reset: boolean := true;
    constant cReset_active_level: std_logic := '0';

end package;
